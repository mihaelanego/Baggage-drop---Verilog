// this module was automatically generated to match the expected results
// for all the possilbe 8-bit numbers

module square_root (
	output reg [15:0] out,
	input  [7:0] in
);

	reg[15:0] roots[255:0];

	initial begin
		roots[8'd0] = 16'b00000000_00000000; // = 0.00 (expected) real: 0.000
		roots[8'd1] = 16'b00000001_00000000; // = 1.00 (expected) real: 1.000
		roots[8'd2] = 16'b00000001_01101010; // = 1.41 (expected) real: 1.414
		roots[8'd3] = 16'b00000001_10111011; // = 1.73 (expected) real: 1.732
		roots[8'd4] = 16'b00000010_00000000; // = 2.00 (expected) real: 2.000
		roots[8'd5] = 16'b00000010_00111100; // = 2.23 (expected) real: 2.236
		roots[8'd6] = 16'b00000010_01110011; // = 2.45 (expected) real: 2.449
		roots[8'd7] = 16'b00000010_10100101; // = 2.64 (expected) real: 2.646
		roots[8'd8] = 16'b00000010_11010100; // = 2.83 (expected) real: 2.828
		roots[8'd9] = 16'b00000011_00000000; // = 3.00 (expected) real: 3.000
		roots[8'd10] = 16'b00000011_00101001; // = 3.16 (expected) real: 3.162
		roots[8'd11] = 16'b00000011_01010001; // = 3.32 (expected) real: 3.317
		roots[8'd12] = 16'b00000011_01110110; // = 3.46 (expected) real: 3.464
		roots[8'd13] = 16'b00000011_10011011; // = 3.61 (expected) real: 3.606
		roots[8'd14] = 16'b00000011_10111101; // = 3.74 (expected) real: 3.742
		roots[8'd15] = 16'b00000011_11011111; // = 3.87 (expected) real: 3.873
		roots[8'd16] = 16'b00000100_00000000; // = 4.00 (expected) real: 4.000
		roots[8'd17] = 16'b00000100_00011111; // = 4.12 (expected) real: 4.123
		roots[8'd18] = 16'b00000100_00111110; // = 4.24 (expected) real: 4.243
		roots[8'd19] = 16'b00000100_01011011; // = 4.36 (expected) real: 4.359
		roots[8'd20] = 16'b00000100_01111000; // = 4.47 (expected) real: 4.472
		roots[8'd21] = 16'b00000100_10010101; // = 4.58 (expected) real: 4.583
		roots[8'd22] = 16'b00000100_10110000; // = 4.69 (expected) real: 4.690
		roots[8'd23] = 16'b00000100_11001011; // = 4.79 (expected) real: 4.796
		roots[8'd24] = 16'b00000100_11100110; // = 4.90 (expected) real: 4.899
		roots[8'd25] = 16'b00000101_00000000; // = 5.00 (expected) real: 5.000
		roots[8'd26] = 16'b00000101_00011001; // = 5.10 (expected) real: 5.099
		roots[8'd27] = 16'b00000101_00110010; // = 5.20 (expected) real: 5.196
		roots[8'd28] = 16'b00000101_01001010; // = 5.29 (expected) real: 5.292
		roots[8'd29] = 16'b00000101_01100010; // = 5.38 (expected) real: 5.385
		roots[8'd30] = 16'b00000101_01111010; // = 5.48 (expected) real: 5.477
		roots[8'd31] = 16'b00000101_10010001; // = 5.57 (expected) real: 5.568
		roots[8'd32] = 16'b00000101_10101000; // = 5.66 (expected) real: 5.657
		roots[8'd33] = 16'b00000101_10111110; // = 5.74 (expected) real: 5.745
		roots[8'd34] = 16'b00000101_11010100; // = 5.83 (expected) real: 5.831
		roots[8'd35] = 16'b00000101_11101010; // = 5.91 (expected) real: 5.916
		roots[8'd36] = 16'b00000110_00000000; // = 6.00 (expected) real: 6.000
		roots[8'd37] = 16'b00000110_00010101; // = 6.08 (expected) real: 6.083
		roots[8'd38] = 16'b00000110_00101010; // = 6.16 (expected) real: 6.164
		roots[8'd39] = 16'b00000110_00111110; // = 6.24 (expected) real: 6.245
		roots[8'd40] = 16'b00000110_01010011; // = 6.32 (expected) real: 6.325
		roots[8'd41] = 16'b00000110_01100111; // = 6.40 (expected) real: 6.403
		roots[8'd42] = 16'b00000110_01111011; // = 6.48 (expected) real: 6.481
		roots[8'd43] = 16'b00000110_10001110; // = 6.55 (expected) real: 6.557
		roots[8'd44] = 16'b00000110_10100010; // = 6.63 (expected) real: 6.633
		roots[8'd45] = 16'b00000110_10110101; // = 6.71 (expected) real: 6.708
		roots[8'd46] = 16'b00000110_11001000; // = 6.78 (expected) real: 6.782
		roots[8'd47] = 16'b00000110_11011011; // = 6.86 (expected) real: 6.856
		roots[8'd48] = 16'b00000110_11101101; // = 6.93 (expected) real: 6.928
		roots[8'd49] = 16'b00000111_00000000; // = 7.00 (expected) real: 7.000
		roots[8'd50] = 16'b00000111_00010010; // = 7.07 (expected) real: 7.071
		roots[8'd51] = 16'b00000111_00100100; // = 7.14 (expected) real: 7.141
		roots[8'd52] = 16'b00000111_00110110; // = 7.21 (expected) real: 7.211
		roots[8'd53] = 16'b00000111_01000111; // = 7.28 (expected) real: 7.280
		roots[8'd54] = 16'b00000111_01011001; // = 7.35 (expected) real: 7.348
		roots[8'd55] = 16'b00000111_01101010; // = 7.41 (expected) real: 7.416
		roots[8'd56] = 16'b00000111_01111011; // = 7.48 (expected) real: 7.483
		roots[8'd57] = 16'b00000111_10001100; // = 7.55 (expected) real: 7.550
		roots[8'd58] = 16'b00000111_10011101; // = 7.61 (expected) real: 7.616
		roots[8'd59] = 16'b00000111_10101110; // = 7.68 (expected) real: 7.681
		roots[8'd60] = 16'b00000111_10111110; // = 7.74 (expected) real: 7.746
		roots[8'd61] = 16'b00000111_11001111; // = 7.81 (expected) real: 7.810
		roots[8'd62] = 16'b00000111_11011111; // = 7.87 (expected) real: 7.874
		roots[8'd63] = 16'b00000111_11101111; // = 7.93 (expected) real: 7.937
		roots[8'd64] = 16'b00001000_00000000; // = 8.00 (expected) real: 8.000
		roots[8'd65] = 16'b00001000_00001111; // = 8.06 (expected) real: 8.062
		roots[8'd66] = 16'b00001000_00011111; // = 8.12 (expected) real: 8.124
		roots[8'd67] = 16'b00001000_00101111; // = 8.18 (expected) real: 8.185
		roots[8'd68] = 16'b00001000_00111111; // = 8.25 (expected) real: 8.246
		roots[8'd69] = 16'b00001000_01001110; // = 8.30 (expected) real: 8.307
		roots[8'd70] = 16'b00001000_01011101; // = 8.36 (expected) real: 8.367
		roots[8'd71] = 16'b00001000_01101101; // = 8.43 (expected) real: 8.426
		roots[8'd72] = 16'b00001000_01111100; // = 8.48 (expected) real: 8.485
		roots[8'd73] = 16'b00001000_10001011; // = 8.54 (expected) real: 8.544
		roots[8'd74] = 16'b00001000_10011010; // = 8.60 (expected) real: 8.602
		roots[8'd75] = 16'b00001000_10101001; // = 8.66 (expected) real: 8.660
		roots[8'd76] = 16'b00001000_10110111; // = 8.71 (expected) real: 8.718
		roots[8'd77] = 16'b00001000_11000110; // = 8.77 (expected) real: 8.775
		roots[8'd78] = 16'b00001000_11010100; // = 8.83 (expected) real: 8.832
		roots[8'd79] = 16'b00001000_11100011; // = 8.89 (expected) real: 8.888
		roots[8'd80] = 16'b00001000_11110001; // = 8.94 (expected) real: 8.944
		roots[8'd81] = 16'b00001001_00000000; // = 9.00 (expected) real: 9.000
		roots[8'd82] = 16'b00001001_00001110; // = 9.05 (expected) real: 9.055
		roots[8'd83] = 16'b00001001_00011100; // = 9.11 (expected) real: 9.110
		roots[8'd84] = 16'b00001001_00101010; // = 9.16 (expected) real: 9.165
		roots[8'd85] = 16'b00001001_00111000; // = 9.22 (expected) real: 9.220
		roots[8'd86] = 16'b00001001_01000110; // = 9.27 (expected) real: 9.274
		roots[8'd87] = 16'b00001001_01010011; // = 9.32 (expected) real: 9.327
		roots[8'd88] = 16'b00001001_01100001; // = 9.38 (expected) real: 9.381
		roots[8'd89] = 16'b00001001_01101111; // = 9.43 (expected) real: 9.434
		roots[8'd90] = 16'b00001001_01111100; // = 9.48 (expected) real: 9.487
		roots[8'd91] = 16'b00001001_10001010; // = 9.54 (expected) real: 9.539
		roots[8'd92] = 16'b00001001_10010111; // = 9.59 (expected) real: 9.592
		roots[8'd93] = 16'b00001001_10100100; // = 9.64 (expected) real: 9.644
		roots[8'd94] = 16'b00001001_10110010; // = 9.70 (expected) real: 9.695
		roots[8'd95] = 16'b00001001_10111111; // = 9.75 (expected) real: 9.747
		roots[8'd96] = 16'b00001001_11001100; // = 9.80 (expected) real: 9.798
		roots[8'd97] = 16'b00001001_11011001; // = 9.85 (expected) real: 9.849
		roots[8'd98] = 16'b00001001_11100110; // = 9.90 (expected) real: 9.899
		roots[8'd99] = 16'b00001001_11110011; // = 9.95 (expected) real: 9.950
		roots[8'd100] = 16'b00001010_00000000; // = 10.00 (expected) real: 10.000
		roots[8'd101] = 16'b00001010_00001100; // = 10.05 (expected) real: 10.050
		roots[8'd102] = 16'b00001010_00011001; // = 10.10 (expected) real: 10.100
		roots[8'd103] = 16'b00001010_00100110; // = 10.15 (expected) real: 10.149
		roots[8'd104] = 16'b00001010_00110010; // = 10.20 (expected) real: 10.198
		roots[8'd105] = 16'b00001010_00111111; // = 10.25 (expected) real: 10.247
		roots[8'd106] = 16'b00001010_01001011; // = 10.29 (expected) real: 10.296
		roots[8'd107] = 16'b00001010_01011000; // = 10.34 (expected) real: 10.344
		roots[8'd108] = 16'b00001010_01100100; // = 10.39 (expected) real: 10.392
		roots[8'd109] = 16'b00001010_01110000; // = 10.44 (expected) real: 10.440
		roots[8'd110] = 16'b00001010_01111100; // = 10.48 (expected) real: 10.488
		roots[8'd111] = 16'b00001010_10001001; // = 10.54 (expected) real: 10.536
		roots[8'd112] = 16'b00001010_10010101; // = 10.58 (expected) real: 10.583
		roots[8'd113] = 16'b00001010_10100001; // = 10.63 (expected) real: 10.630
		roots[8'd114] = 16'b00001010_10101101; // = 10.68 (expected) real: 10.677
		roots[8'd115] = 16'b00001010_10111001; // = 10.72 (expected) real: 10.724
		roots[8'd116] = 16'b00001010_11000101; // = 10.77 (expected) real: 10.770
		roots[8'd117] = 16'b00001010_11010001; // = 10.82 (expected) real: 10.817
		roots[8'd118] = 16'b00001010_11011100; // = 10.86 (expected) real: 10.863
		roots[8'd119] = 16'b00001010_11101000; // = 10.91 (expected) real: 10.909
		roots[8'd120] = 16'b00001010_11110100; // = 10.95 (expected) real: 10.954
		roots[8'd121] = 16'b00001011_00000000; // = 11.00 (expected) real: 11.000
		roots[8'd122] = 16'b00001011_00001011; // = 11.04 (expected) real: 11.045
		roots[8'd123] = 16'b00001011_00010111; // = 11.09 (expected) real: 11.091
		roots[8'd124] = 16'b00001011_00100010; // = 11.13 (expected) real: 11.136
		roots[8'd125] = 16'b00001011_00101110; // = 11.18 (expected) real: 11.180
		roots[8'd126] = 16'b00001011_00111001; // = 11.22 (expected) real: 11.225
		roots[8'd127] = 16'b00001011_01000100; // = 11.27 (expected) real: 11.269
		roots[8'd128] = 16'b00001011_01010000; // = 11.31 (expected) real: 11.314
		roots[8'd129] = 16'b00001011_01011011; // = 11.36 (expected) real: 11.358
		roots[8'd130] = 16'b00001011_01100110; // = 11.40 (expected) real: 11.402
		roots[8'd131] = 16'b00001011_01110010; // = 11.45 (expected) real: 11.446
		roots[8'd132] = 16'b00001011_01111101; // = 11.49 (expected) real: 11.489
		roots[8'd133] = 16'b00001011_10001000; // = 11.53 (expected) real: 11.533
		roots[8'd134] = 16'b00001011_10010011; // = 11.57 (expected) real: 11.576
		roots[8'd135] = 16'b00001011_10011110; // = 11.62 (expected) real: 11.619
		roots[8'd136] = 16'b00001011_10101001; // = 11.66 (expected) real: 11.662
		roots[8'd137] = 16'b00001011_10110100; // = 11.70 (expected) real: 11.705
		roots[8'd138] = 16'b00001011_10111111; // = 11.75 (expected) real: 11.747
		roots[8'd139] = 16'b00001011_11001010; // = 11.79 (expected) real: 11.790
		roots[8'd140] = 16'b00001011_11010101; // = 11.83 (expected) real: 11.832
		roots[8'd141] = 16'b00001011_11011111; // = 11.87 (expected) real: 11.874
		roots[8'd142] = 16'b00001011_11101010; // = 11.91 (expected) real: 11.916
		roots[8'd143] = 16'b00001011_11110101; // = 11.96 (expected) real: 11.958
		roots[8'd144] = 16'b00001100_00000000; // = 12.00 (expected) real: 12.000
		roots[8'd145] = 16'b00001100_00001010; // = 12.04 (expected) real: 12.042
		roots[8'd146] = 16'b00001100_00010101; // = 12.08 (expected) real: 12.083
		roots[8'd147] = 16'b00001100_00011111; // = 12.12 (expected) real: 12.124
		roots[8'd148] = 16'b00001100_00101010; // = 12.16 (expected) real: 12.166
		roots[8'd149] = 16'b00001100_00110100; // = 12.20 (expected) real: 12.207
		roots[8'd150] = 16'b00001100_00111111; // = 12.25 (expected) real: 12.247
		roots[8'd151] = 16'b00001100_01001001; // = 12.29 (expected) real: 12.288
		roots[8'd152] = 16'b00001100_01010100; // = 12.33 (expected) real: 12.329
		roots[8'd153] = 16'b00001100_01011110; // = 12.37 (expected) real: 12.369
		roots[8'd154] = 16'b00001100_01101000; // = 12.41 (expected) real: 12.410
		roots[8'd155] = 16'b00001100_01110011; // = 12.45 (expected) real: 12.450
		roots[8'd156] = 16'b00001100_01111101; // = 12.49 (expected) real: 12.490
		roots[8'd157] = 16'b00001100_10000111; // = 12.53 (expected) real: 12.530
		roots[8'd158] = 16'b00001100_10010001; // = 12.57 (expected) real: 12.570
		roots[8'd159] = 16'b00001100_10011100; // = 12.61 (expected) real: 12.610
		roots[8'd160] = 16'b00001100_10100110; // = 12.65 (expected) real: 12.649
		roots[8'd161] = 16'b00001100_10110000; // = 12.69 (expected) real: 12.689
		roots[8'd162] = 16'b00001100_10111010; // = 12.73 (expected) real: 12.728
		roots[8'd163] = 16'b00001100_11000100; // = 12.77 (expected) real: 12.767
		roots[8'd164] = 16'b00001100_11001110; // = 12.80 (expected) real: 12.806
		roots[8'd165] = 16'b00001100_11011000; // = 12.84 (expected) real: 12.845
		roots[8'd166] = 16'b00001100_11100010; // = 12.88 (expected) real: 12.884
		roots[8'd167] = 16'b00001100_11101100; // = 12.92 (expected) real: 12.923
		roots[8'd168] = 16'b00001100_11110110; // = 12.96 (expected) real: 12.961
		roots[8'd169] = 16'b00001101_00000000; // = 13.00 (expected) real: 13.000
		roots[8'd170] = 16'b00001101_00001001; // = 13.04 (expected) real: 13.038
		roots[8'd171] = 16'b00001101_00010011; // = 13.07 (expected) real: 13.077
		roots[8'd172] = 16'b00001101_00011101; // = 13.11 (expected) real: 13.115
		roots[8'd173] = 16'b00001101_00100111; // = 13.15 (expected) real: 13.153
		roots[8'd174] = 16'b00001101_00110000; // = 13.19 (expected) real: 13.191
		roots[8'd175] = 16'b00001101_00111010; // = 13.23 (expected) real: 13.229
		roots[8'd176] = 16'b00001101_01000100; // = 13.27 (expected) real: 13.266
		roots[8'd177] = 16'b00001101_01001101; // = 13.30 (expected) real: 13.304
		roots[8'd178] = 16'b00001101_01010111; // = 13.34 (expected) real: 13.342
		roots[8'd179] = 16'b00001101_01100001; // = 13.38 (expected) real: 13.379
		roots[8'd180] = 16'b00001101_01101010; // = 13.41 (expected) real: 13.416
		roots[8'd181] = 16'b00001101_01110100; // = 13.45 (expected) real: 13.454
		roots[8'd182] = 16'b00001101_01111101; // = 13.49 (expected) real: 13.491
		roots[8'd183] = 16'b00001101_10000111; // = 13.53 (expected) real: 13.528
		roots[8'd184] = 16'b00001101_10010000; // = 13.56 (expected) real: 13.565
		roots[8'd185] = 16'b00001101_10011001; // = 13.60 (expected) real: 13.601
		roots[8'd186] = 16'b00001101_10100011; // = 13.64 (expected) real: 13.638
		roots[8'd187] = 16'b00001101_10101100; // = 13.67 (expected) real: 13.675
		roots[8'd188] = 16'b00001101_10110110; // = 13.71 (expected) real: 13.711
		roots[8'd189] = 16'b00001101_10111111; // = 13.75 (expected) real: 13.748
		roots[8'd190] = 16'b00001101_11001000; // = 13.78 (expected) real: 13.784
		roots[8'd191] = 16'b00001101_11010001; // = 13.82 (expected) real: 13.820
		roots[8'd192] = 16'b00001101_11011011; // = 13.86 (expected) real: 13.856
		roots[8'd193] = 16'b00001101_11100100; // = 13.89 (expected) real: 13.892
		roots[8'd194] = 16'b00001101_11101101; // = 13.93 (expected) real: 13.928
		roots[8'd195] = 16'b00001101_11110110; // = 13.96 (expected) real: 13.964
		roots[8'd196] = 16'b00001110_00000000; // = 14.00 (expected) real: 14.000
		roots[8'd197] = 16'b00001110_00001001; // = 14.04 (expected) real: 14.036
		roots[8'd198] = 16'b00001110_00010010; // = 14.07 (expected) real: 14.071
		roots[8'd199] = 16'b00001110_00011011; // = 14.11 (expected) real: 14.107
		roots[8'd200] = 16'b00001110_00100100; // = 14.14 (expected) real: 14.142
		roots[8'd201] = 16'b00001110_00101101; // = 14.18 (expected) real: 14.177
		roots[8'd202] = 16'b00001110_00110110; // = 14.21 (expected) real: 14.213
		roots[8'd203] = 16'b00001110_00111111; // = 14.25 (expected) real: 14.248
		roots[8'd204] = 16'b00001110_01001000; // = 14.28 (expected) real: 14.283
		roots[8'd205] = 16'b00001110_01010001; // = 14.32 (expected) real: 14.318
		roots[8'd206] = 16'b00001110_01011010; // = 14.35 (expected) real: 14.353
		roots[8'd207] = 16'b00001110_01100011; // = 14.39 (expected) real: 14.387
		roots[8'd208] = 16'b00001110_01101100; // = 14.42 (expected) real: 14.422
		roots[8'd209] = 16'b00001110_01110100; // = 14.45 (expected) real: 14.457
		roots[8'd210] = 16'b00001110_01111101; // = 14.49 (expected) real: 14.491
		roots[8'd211] = 16'b00001110_10000110; // = 14.52 (expected) real: 14.526
		roots[8'd212] = 16'b00001110_10001111; // = 14.56 (expected) real: 14.560
		roots[8'd213] = 16'b00001110_10011000; // = 14.59 (expected) real: 14.595
		roots[8'd214] = 16'b00001110_10100000; // = 14.63 (expected) real: 14.629
		roots[8'd215] = 16'b00001110_10101001; // = 14.66 (expected) real: 14.663
		roots[8'd216] = 16'b00001110_10110010; // = 14.70 (expected) real: 14.697
		roots[8'd217] = 16'b00001110_10111011; // = 14.73 (expected) real: 14.731
		roots[8'd218] = 16'b00001110_11000011; // = 14.76 (expected) real: 14.765
		roots[8'd219] = 16'b00001110_11001100; // = 14.80 (expected) real: 14.799
		roots[8'd220] = 16'b00001110_11010101; // = 14.83 (expected) real: 14.832
		roots[8'd221] = 16'b00001110_11011101; // = 14.86 (expected) real: 14.866
		roots[8'd222] = 16'b00001110_11100110; // = 14.90 (expected) real: 14.900
		roots[8'd223] = 16'b00001110_11101110; // = 14.93 (expected) real: 14.933
		roots[8'd224] = 16'b00001110_11110111; // = 14.96 (expected) real: 14.967
		roots[8'd225] = 16'b00001111_00000000; // = 15.00 (expected) real: 15.000
		roots[8'd226] = 16'b00001111_00001000; // = 15.03 (expected) real: 15.033
		roots[8'd227] = 16'b00001111_00010001; // = 15.07 (expected) real: 15.067
		roots[8'd228] = 16'b00001111_00011001; // = 15.10 (expected) real: 15.100
		roots[8'd229] = 16'b00001111_00100001; // = 15.13 (expected) real: 15.133
		roots[8'd230] = 16'b00001111_00101010; // = 15.16 (expected) real: 15.166
		roots[8'd231] = 16'b00001111_00110010; // = 15.20 (expected) real: 15.199
		roots[8'd232] = 16'b00001111_00111011; // = 15.23 (expected) real: 15.232
		roots[8'd233] = 16'b00001111_01000011; // = 15.26 (expected) real: 15.264
		roots[8'd234] = 16'b00001111_01001100; // = 15.30 (expected) real: 15.297
		roots[8'd235] = 16'b00001111_01010100; // = 15.33 (expected) real: 15.330
		roots[8'd236] = 16'b00001111_01011100; // = 15.36 (expected) real: 15.362
		roots[8'd237] = 16'b00001111_01100101; // = 15.39 (expected) real: 15.395
		roots[8'd238] = 16'b00001111_01101101; // = 15.43 (expected) real: 15.427
		roots[8'd239] = 16'b00001111_01110101; // = 15.46 (expected) real: 15.460
		roots[8'd240] = 16'b00001111_01111101; // = 15.49 (expected) real: 15.492
		roots[8'd241] = 16'b00001111_10000110; // = 15.52 (expected) real: 15.524
		roots[8'd242] = 16'b00001111_10001110; // = 15.55 (expected) real: 15.556
		roots[8'd243] = 16'b00001111_10010110; // = 15.59 (expected) real: 15.588
		roots[8'd244] = 16'b00001111_10011110; // = 15.62 (expected) real: 15.620
		roots[8'd245] = 16'b00001111_10100111; // = 15.65 (expected) real: 15.652
		roots[8'd246] = 16'b00001111_10101111; // = 15.68 (expected) real: 15.684
		roots[8'd247] = 16'b00001111_10110111; // = 15.71 (expected) real: 15.716
		roots[8'd248] = 16'b00001111_10111111; // = 15.75 (expected) real: 15.748
		roots[8'd249] = 16'b00001111_11000111; // = 15.78 (expected) real: 15.780
		roots[8'd250] = 16'b00001111_11001111; // = 15.81 (expected) real: 15.811
		roots[8'd251] = 16'b00001111_11010111; // = 15.84 (expected) real: 15.843
		roots[8'd252] = 16'b00001111_11011111; // = 15.87 (expected) real: 15.875
		roots[8'd253] = 16'b00001111_11100111; // = 15.90 (expected) real: 15.906
		roots[8'd254] = 16'b00001111_11101111; // = 15.93 (expected) real: 15.937
		roots[8'd255] = 16'b00001111_11110111; // = 15.96 (expected) real: 15.969
	end

	always @(in) begin
		out = roots[in];
	end
endmodule